let gmbs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[gm]
let gds_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[vth]
let id_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[id]
let ibd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[gbs]
let isub_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[isub]
let igidl_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[igisl]
let igs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[igs]
let igd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[igd]
let igb_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[igb]
let igcs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[vgs]
let vds_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[vds]
let cgg_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cdd]
let cds_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cds]
let csg_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[csg]
let csd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[csd]
let css_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[css]
let cgb_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cdb]
let csb_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[csb]
let cbb_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M0=@m.x1.XM0.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[gm]
let gds_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[vth]
let id_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[id]
let ibd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[gbs]
let isub_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[isub]
let igidl_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[igisl]
let igs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[igs]
let igd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[igd]
let igb_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[igb]
let igcs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[vgs]
let vds_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[vds]
let cgg_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cdd]
let cds_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cds]
let csg_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[csg]
let csd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[csd]
let css_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[css]
let cgb_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cdb]
let csb_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[csb]
let cbb_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M1=@m.x1.XM1.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[gm]
let gds_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[vth]
let id_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[id]
let ibd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[gbs]
let isub_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[isub]
let igidl_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[igisl]
let igs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[igs]
let igd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[igd]
let igb_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[igb]
let igcs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[vgs]
let vds_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[vds]
let cgg_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cdd]
let cds_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cds]
let csg_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[csg]
let csd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[csd]
let css_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[css]
let cgb_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cdb]
let csb_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[csb]
let cbb_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M2=@m.x1.XM2.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[gm]
let gds_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[vth]
let id_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[id]
let ibd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[gbs]
let isub_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[isub]
let igidl_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[igisl]
let igs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[igs]
let igd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[igd]
let igb_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[igb]
let igcs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[vgs]
let vds_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[vds]
let cgg_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cdd]
let cds_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cds]
let csg_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[csg]
let csd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[csd]
let css_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[css]
let cgb_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cdb]
let csb_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[csb]
let cbb_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M3=@m.x1.XM3.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[gm]
let gds_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[vth]
let id_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[id]
let ibd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[gbs]
let isub_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[isub]
let igidl_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[igisl]
let igs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[igs]
let igd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[igd]
let igb_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[igb]
let igcs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[vgs]
let vds_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[vds]
let cgg_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cdd]
let cds_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cds]
let csg_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[csg]
let csd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[csd]
let css_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[css]
let cgb_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cdb]
let csb_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[csb]
let cbb_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M4=@m.x1.XM4.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[gm]
let gds_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[vth]
let id_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[id]
let ibd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[gbs]
let isub_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[isub]
let igidl_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[igisl]
let igs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[igs]
let igd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[igd]
let igb_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[igb]
let igcs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[vgs]
let vds_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[vds]
let cgg_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cdd]
let cds_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cds]
let csg_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[csg]
let csd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[csd]
let css_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[css]
let cgb_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cdb]
let csb_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[csb]
let cbb_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M5=@m.x1.XM5.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[gm]
let gds_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[vth]
let id_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[id]
let ibd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[gbs]
let isub_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[isub]
let igidl_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[igisl]
let igs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[igs]
let igd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[igd]
let igb_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[igb]
let igcs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[vgs]
let vds_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[vds]
let cgg_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cdd]
let cds_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cds]
let csg_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[csg]
let csd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[csd]
let css_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[css]
let cgb_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cdb]
let csb_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[csb]
let cbb_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M6=@m.x1.XM6.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[gm]
let gds_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[vth]
let id_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[id]
let ibd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[gbs]
let isub_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[isub]
let igidl_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[igisl]
let igs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[igs]
let igd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[igd]
let igb_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[igb]
let igcs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[vgs]
let vds_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[vds]
let cgg_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cdd]
let cds_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cds]
let csg_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[csg]
let csd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[csd]
let css_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[css]
let cgb_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cdb]
let csb_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[csb]
let cbb_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M7=@m.x1.XM7.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[gm]
let gds_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[vth]
let id_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[id]
let ibd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[gbs]
let isub_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[isub]
let igidl_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[igisl]
let igs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[igs]
let igd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[igd]
let igb_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[igb]
let igcs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[vgs]
let vds_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[vds]
let cgg_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cdd]
let cds_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cds]
let csg_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[csg]
let csd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[csd]
let css_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[css]
let cgb_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cdb]
let csb_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[csb]
let cbb_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M8=@m.x1.XM8.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[gm]
let gds_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[vth]
let id_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[id]
let ibd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[gbs]
let isub_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[isub]
let igidl_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[igisl]
let igs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[igs]
let igd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[igd]
let igb_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[igb]
let igcs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[vgs]
let vds_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[vds]
let cgg_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cdd]
let cds_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cds]
let csg_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[csg]
let csd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[csd]
let css_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[css]
let cgb_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cdb]
let csb_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[csb]
let cbb_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M9=@m.x1.XM9.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[gm]
let gds_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[vth]
let id_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[id]
let ibd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[gbs]
let isub_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[isub]
let igidl_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[igisl]
let igs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[igs]
let igd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[igd]
let igb_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[igb]
let igcs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[vgs]
let vds_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[vds]
let cgg_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cdd]
let cds_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cds]
let csg_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[csg]
let csd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[csd]
let css_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[css]
let cgb_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cdb]
let csb_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[csb]
let cbb_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M10=@m.x1.XM10.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[gmbs]
let gm_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[gm]
let gds_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[gds]
let vdsat_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[vdsat]
let vth_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[vth]
let id_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[id]
let ibd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[ibd]
let ibs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[ibs]
let gbd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[gbd]
let gbs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[gbs]
let isub_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[isub]
let igidl_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[igidl]
let igisl_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[igisl]
let igs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[igs]
let igd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[igd]
let igb_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[igb]
let igcs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[igcs]
let vbs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[vbs]
let vgs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[vgs]
let vds_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[vds]
let cgg_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cgg]
let cgs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cgs]
let cgd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cgd]
let cbg_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cbg]
let cbd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cbd]
let cbs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cbs]
let cdg_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cdg]
let cdd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cdd]
let cds_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cds]
let csg_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[csg]
let csd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[csd]
let css_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[css]
let cgb_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cgb]
let cdb_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cdb]
let csb_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[csb]
let cbb_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[cbb]
let capbd_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[capbd]
let capbs_M11=@m.x1.XM11.msky130_fd_pr__pfet_01v8[capbs]

let gmbs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[gm]
let gds_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[vth]
let id_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[id]
let ibd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[gbs]
let isub_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[isub]
let igidl_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[igisl]
let igs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[igs]
let igd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[igd]
let igb_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[igb]
let igcs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[vgs]
let vds_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[vds]
let cgg_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cdd]
let cds_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cds]
let csg_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[csg]
let csd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[csd]
let css_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[css]
let cgb_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cdb]
let csb_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[csb]
let cbb_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M12=@m.x1.XM12.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[gm]
let gds_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[vth]
let id_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[id]
let ibd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[gbs]
let isub_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[isub]
let igidl_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[igisl]
let igs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[igs]
let igd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[igd]
let igb_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[igb]
let igcs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[vgs]
let vds_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[vds]
let cgg_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cdd]
let cds_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cds]
let csg_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[csg]
let csd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[csd]
let css_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[css]
let cgb_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cdb]
let csb_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[csb]
let cbb_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M13=@m.x1.XM13.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[gm]
let gds_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[vth]
let id_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[id]
let ibd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[gbs]
let isub_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[isub]
let igidl_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[igisl]
let igs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[igs]
let igd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[igd]
let igb_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[igb]
let igcs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[vgs]
let vds_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[vds]
let cgg_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cdd]
let cds_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cds]
let csg_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[csg]
let csd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[csd]
let css_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[css]
let cgb_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cdb]
let csb_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[csb]
let cbb_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M14=@m.x1.XM14.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[gm]
let gds_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[vth]
let id_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[id]
let ibd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[gbs]
let isub_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[isub]
let igidl_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[igisl]
let igs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[igs]
let igd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[igd]
let igb_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[igb]
let igcs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[vgs]
let vds_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[vds]
let cgg_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cdd]
let cds_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cds]
let csg_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[csg]
let csd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[csd]
let css_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[css]
let cgb_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cdb]
let csb_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[csb]
let cbb_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M15=@m.x1.XM15.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[gm]
let gds_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[vth]
let id_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[id]
let ibd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[gbs]
let isub_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[isub]
let igidl_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[igisl]
let igs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[igs]
let igd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[igd]
let igb_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[igb]
let igcs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[vgs]
let vds_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[vds]
let cgg_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cdd]
let cds_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cds]
let csg_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[csg]
let csd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[csd]
let css_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[css]
let cgb_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cdb]
let csb_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[csb]
let cbb_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M16=@m.x1.XM16.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[gm]
let gds_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[vth]
let id_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[id]
let ibd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[gbs]
let isub_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[isub]
let igidl_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[igisl]
let igs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[igs]
let igd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[igd]
let igb_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[igb]
let igcs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[vgs]
let vds_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[vds]
let cgg_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cdd]
let cds_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cds]
let csg_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[csg]
let csd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[csd]
let css_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[css]
let cgb_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cdb]
let csb_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[csb]
let cbb_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M17=@m.x1.XM17.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[gm]
let gds_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[vth]
let id_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[id]
let ibd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[gbs]
let isub_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[isub]
let igidl_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[igisl]
let igs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[igs]
let igd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[igd]
let igb_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[igb]
let igcs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[vgs]
let vds_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[vds]
let cgg_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cdd]
let cds_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cds]
let csg_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[csg]
let csd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[csd]
let css_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[css]
let cgb_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cdb]
let csb_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[csb]
let cbb_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M18=@m.x1.XM18.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[gm]
let gds_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[vth]
let id_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[id]
let ibd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[gbs]
let isub_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[isub]
let igidl_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[igisl]
let igs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[igs]
let igd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[igd]
let igb_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[igb]
let igcs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[vgs]
let vds_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[vds]
let cgg_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cdd]
let cds_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cds]
let csg_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[csg]
let csd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[csd]
let css_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[css]
let cgb_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cdb]
let csb_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[csb]
let cbb_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M19=@m.x1.XM19.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[gm]
let gds_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[vth]
let id_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[id]
let ibd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[gbs]
let isub_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[isub]
let igidl_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[igisl]
let igs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[igs]
let igd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[igd]
let igb_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[igb]
let igcs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[vgs]
let vds_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[vds]
let cgg_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cdd]
let cds_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cds]
let csg_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[csg]
let csd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[csd]
let css_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[css]
let cgb_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cdb]
let csb_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[csb]
let cbb_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M20=@m.x1.XM20.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[gm]
let gds_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[vth]
let id_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[id]
let ibd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[gbs]
let isub_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[isub]
let igidl_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[igisl]
let igs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[igs]
let igd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[igd]
let igb_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[igb]
let igcs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[vgs]
let vds_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[vds]
let cgg_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cdd]
let cds_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cds]
let csg_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[csg]
let csd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[csd]
let css_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[css]
let cgb_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cdb]
let csb_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[csb]
let cbb_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M21=@m.x1.XM21.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[gm]
let gds_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[vth]
let id_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[id]
let ibd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[gbs]
let isub_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[isub]
let igidl_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[igisl]
let igs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[igs]
let igd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[igd]
let igb_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[igb]
let igcs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[vgs]
let vds_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[vds]
let cgg_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cdd]
let cds_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cds]
let csg_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[csg]
let csd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[csd]
let css_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[css]
let cgb_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cdb]
let csb_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[csb]
let cbb_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M22=@m.x1.XM22.msky130_fd_pr__nfet_01v8[capbs]

let gmbs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[gmbs]
let gm_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[gm]
let gds_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[gds]
let vdsat_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[vdsat]
let vth_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[vth]
let id_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[id]
let ibd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[ibd]
let ibs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[ibs]
let gbd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[gbd]
let gbs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[gbs]
let isub_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[isub]
let igidl_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[igidl]
let igisl_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[igisl]
let igs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[igs]
let igd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[igd]
let igb_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[igb]
let igcs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[igcs]
let vbs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[vbs]
let vgs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[vgs]
let vds_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[vds]
let cgg_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cgg]
let cgs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cgs]
let cgd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cgd]
let cbg_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cbg]
let cbd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cbd]
let cbs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cbs]
let cdg_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cdg]
let cdd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cdd]
let cds_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cds]
let csg_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[csg]
let csd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[csd]
let css_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[css]
let cgb_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cgb]
let cdb_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cdb]
let csb_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[csb]
let cbb_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[cbb]
let capbd_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[capbd]
let capbs_M23=@m.x1.XM23.msky130_fd_pr__nfet_01v8[capbs]

let dc_Ib=@Ib[dc]
let acmag_Ib=@Ib[acmag]
let acphase_Ib=@Ib[acphase]
let acreal_Ib=@Ib[acreal]
let acimag_Ib=@Ib[acimag]
let v_Ib=@Ib[v]
let p_Ib=@Ib[p]
let current_Ib=@Ib[current]

let capacitance_C0=@c.x1.XC0.c1[capacitance]
let cap_C0=@c.x1.XC0.c1[cap]
let c_C0=@c.x1.XC0.c1[c]
let ic_C0=@c.x1.XC0.c1[ic]
let temp_C0=@c.x1.XC0.c1[temp]
let dtemp_C0=@c.x1.XC0.c1[dtemp]
let w_C0=@c.x1.XC0.c1[w]
let l_C0=@c.x1.XC0.c1[l]
let m_C0=@c.x1.XC0.c1[m]
let scale_C0=@c.x1.XC0.c1[scale]
let i_C0=@c.x1.XC0.c1[i]
let p_C0=@c.x1.XC0.c1[p]
let sens_dc_C0=@c.x1.XC0.c1[sens_dc]
let sens_real_C0=@c.x1.XC0.c1[sens_real]
let sens_imag_C0=@c.x1.XC0.c1[sens_imag]
let sens_mag_C0=@c.x1.XC0.c1[sens_mag]
let sens_ph_C0=@c.x1.XC0.c1[sens_ph]
let sens_cplx_C0=@c.x1.XC0.c1[sens_cplx]

let capacitance_C1=@c.x1.XC1.c1[capacitance]
let cap_C1=@c.x1.XC1.c1[cap]
let c_C1=@c.x1.XC1.c1[c]
let ic_C1=@c.x1.XC1.c1[ic]
let temp_C1=@c.x1.XC1.c1[temp]
let dtemp_C1=@c.x1.XC1.c1[dtemp]
let w_C1=@c.x1.XC1.c1[w]
let l_C1=@c.x1.XC1.c1[l]
let m_C1=@c.x1.XC1.c1[m]
let scale_C1=@c.x1.XC1.c1[scale]
let i_C1=@c.x1.XC1.c1[i]
let p_C1=@c.x1.XC1.c1[p]
let sens_dc_C1=@c.x1.XC1.c1[sens_dc]
let sens_real_C1=@c.x1.XC1.c1[sens_real]
let sens_imag_C1=@c.x1.XC1.c1[sens_imag]
let sens_mag_C1=@c.x1.XC1.c1[sens_mag]
let sens_ph_C1=@c.x1.XC1.c1[sens_ph]
let sens_cplx_C1=@c.x1.XC1.c1[sens_cplx]

write AMP_NMCF_op gmbs_M0 gm_M0 gds_M0 vdsat_M0 vth_M0 id_M0 ibd_M0 ibs_M0 gbd_M0 gbs_M0 isub_M0 igidl_M0 igisl_M0 igs_M0 igd_M0 igb_M0 igcs_M0 vbs_M0 vgs_M0 vds_M0 cgg_M0 cgs_M0 cgd_M0 cbg_M0 cbd_M0 cbs_M0 cdg_M0 cdd_M0 cds_M0 csg_M0 csd_M0 css_M0 cgb_M0 cdb_M0 csb_M0 cbb_M0 capbd_M0 capbs_M0 gmbs_M1 gm_M1 gds_M1 vdsat_M1 vth_M1 id_M1 ibd_M1 ibs_M1 gbd_M1 gbs_M1 isub_M1 igidl_M1 igisl_M1 igs_M1 igd_M1 igb_M1 igcs_M1 vbs_M1 vgs_M1 vds_M1 cgg_M1 cgs_M1 cgd_M1 cbg_M1 cbd_M1 cbs_M1 cdg_M1 cdd_M1 cds_M1 csg_M1 csd_M1 css_M1 cgb_M1 cdb_M1 csb_M1 cbb_M1 capbd_M1 capbs_M1 gmbs_M2 gm_M2 gds_M2 vdsat_M2 vth_M2 id_M2 ibd_M2 ibs_M2 gbd_M2 gbs_M2 isub_M2 igidl_M2 igisl_M2 igs_M2 igd_M2 igb_M2 igcs_M2 vbs_M2 vgs_M2 vds_M2 cgg_M2 cgs_M2 cgd_M2 cbg_M2 cbd_M2 cbs_M2 cdg_M2 cdd_M2 cds_M2 csg_M2 csd_M2 css_M2 cgb_M2 cdb_M2 csb_M2 cbb_M2 capbd_M2 capbs_M2 gmbs_M3 gm_M3 gds_M3 vdsat_M3 vth_M3 id_M3 ibd_M3 ibs_M3 gbd_M3 gbs_M3 isub_M3 igidl_M3 igisl_M3 igs_M3 igd_M3 igb_M3 igcs_M3 vbs_M3 vgs_M3 vds_M3 cgg_M3 cgs_M3 cgd_M3 cbg_M3 cbd_M3 cbs_M3 cdg_M3 cdd_M3 cds_M3 csg_M3 csd_M3 css_M3 cgb_M3 cdb_M3 csb_M3 cbb_M3 capbd_M3 capbs_M3 gmbs_M4 gm_M4 gds_M4 vdsat_M4 vth_M4 id_M4 ibd_M4 ibs_M4 gbd_M4 gbs_M4 isub_M4 igidl_M4 igisl_M4 igs_M4 igd_M4 igb_M4 igcs_M4 vbs_M4 vgs_M4 vds_M4 cgg_M4 cgs_M4 cgd_M4 cbg_M4 cbd_M4 cbs_M4 cdg_M4 cdd_M4 cds_M4 csg_M4 csd_M4 css_M4 cgb_M4 cdb_M4 csb_M4 cbb_M4 capbd_M4 capbs_M4 gmbs_M5 gm_M5 gds_M5 vdsat_M5 vth_M5 id_M5 ibd_M5 ibs_M5 gbd_M5 gbs_M5 isub_M5 igidl_M5 igisl_M5 igs_M5 igd_M5 igb_M5 igcs_M5 vbs_M5 vgs_M5 vds_M5 cgg_M5 cgs_M5 cgd_M5 cbg_M5 cbd_M5 cbs_M5 cdg_M5 cdd_M5 cds_M5 csg_M5 csd_M5 css_M5 cgb_M5 cdb_M5 csb_M5 cbb_M5 capbd_M5 capbs_M5 gmbs_M6 gm_M6 gds_M6 vdsat_M6 vth_M6 id_M6 ibd_M6 ibs_M6 gbd_M6 gbs_M6 isub_M6 igidl_M6 igisl_M6 igs_M6 igd_M6 igb_M6 igcs_M6 vbs_M6 vgs_M6 vds_M6 cgg_M6 cgs_M6 cgd_M6 cbg_M6 cbd_M6 cbs_M6 cdg_M6 cdd_M6 cds_M6 csg_M6 csd_M6 css_M6 cgb_M6 cdb_M6 csb_M6 cbb_M6 capbd_M6 capbs_M6 gmbs_M7 gm_M7 gds_M7 vdsat_M7 vth_M7 id_M7 ibd_M7 ibs_M7 gbd_M7 gbs_M7 isub_M7 igidl_M7 igisl_M7 igs_M7 igd_M7 igb_M7 igcs_M7 vbs_M7 vgs_M7 vds_M7 cgg_M7 cgs_M7 cgd_M7 cbg_M7 cbd_M7 cbs_M7 cdg_M7 cdd_M7 cds_M7 csg_M7 csd_M7 css_M7 cgb_M7 cdb_M7 csb_M7 cbb_M7 capbd_M7 capbs_M7 gmbs_M8 gm_M8 gds_M8 vdsat_M8 vth_M8 id_M8 ibd_M8 ibs_M8 gbd_M8 gbs_M8 isub_M8 igidl_M8 igisl_M8 igs_M8 igd_M8 igb_M8 igcs_M8 vbs_M8 vgs_M8 vds_M8 cgg_M8 cgs_M8 cgd_M8 cbg_M8 cbd_M8 cbs_M8 cdg_M8 cdd_M8 cds_M8 csg_M8 csd_M8 css_M8 cgb_M8 cdb_M8 csb_M8 cbb_M8 capbd_M8 capbs_M8 gmbs_M9 gm_M9 gds_M9 vdsat_M9 vth_M9 id_M9 ibd_M9 ibs_M9 gbd_M9 gbs_M9 isub_M9 igidl_M9 igisl_M9 igs_M9 igd_M9 igb_M9 igcs_M9 vbs_M9 vgs_M9 vds_M9 cgg_M9 cgs_M9 cgd_M9 cbg_M9 cbd_M9 cbs_M9 cdg_M9 cdd_M9 cds_M9 csg_M9 csd_M9 css_M9 cgb_M9 cdb_M9 csb_M9 cbb_M9 capbd_M9 capbs_M9 gmbs_M10 gm_M10 gds_M10 vdsat_M10 vth_M10 id_M10 ibd_M10 ibs_M10 gbd_M10 gbs_M10 isub_M10 igidl_M10 igisl_M10 igs_M10 igd_M10 igb_M10 igcs_M10 vbs_M10 vgs_M10 vds_M10 cgg_M10 cgs_M10 cgd_M10 cbg_M10 cbd_M10 cbs_M10 cdg_M10 cdd_M10 cds_M10 csg_M10 csd_M10 css_M10 cgb_M10 cdb_M10 csb_M10 cbb_M10 capbd_M10 capbs_M10 gmbs_M11 gm_M11 gds_M11 vdsat_M11 vth_M11 id_M11 ibd_M11 ibs_M11 gbd_M11 gbs_M11 isub_M11 igidl_M11 igisl_M11 igs_M11 igd_M11 igb_M11 igcs_M11 vbs_M11 vgs_M11 vds_M11 cgg_M11 cgs_M11 cgd_M11 cbg_M11 cbd_M11 cbs_M11 cdg_M11 cdd_M11 cds_M11 csg_M11 csd_M11 css_M11 cgb_M11 cdb_M11 csb_M11 cbb_M11 capbd_M11 capbs_M11 gmbs_M12 gm_M12 gds_M12 vdsat_M12 vth_M12 id_M12 ibd_M12 ibs_M12 gbd_M12 gbs_M12 isub_M12 igidl_M12 igisl_M12 igs_M12 igd_M12 igb_M12 igcs_M12 vbs_M12 vgs_M12 vds_M12 cgg_M12 cgs_M12 cgd_M12 cbg_M12 cbd_M12 cbs_M12 cdg_M12 cdd_M12 cds_M12 csg_M12 csd_M12 css_M12 cgb_M12 cdb_M12 csb_M12 cbb_M12 capbd_M12 capbs_M12 gmbs_M13 gm_M13 gds_M13 vdsat_M13 vth_M13 id_M13 ibd_M13 ibs_M13 gbd_M13 gbs_M13 isub_M13 igidl_M13 igisl_M13 igs_M13 igd_M13 igb_M13 igcs_M13 vbs_M13 vgs_M13 vds_M13 cgg_M13 cgs_M13 cgd_M13 cbg_M13 cbd_M13 cbs_M13 cdg_M13 cdd_M13 cds_M13 csg_M13 csd_M13 css_M13 cgb_M13 cdb_M13 csb_M13 cbb_M13 capbd_M13 capbs_M13 gmbs_M14 gm_M14 gds_M14 vdsat_M14 vth_M14 id_M14 ibd_M14 ibs_M14 gbd_M14 gbs_M14 isub_M14 igidl_M14 igisl_M14 igs_M14 igd_M14 igb_M14 igcs_M14 vbs_M14 vgs_M14 vds_M14 cgg_M14 cgs_M14 cgd_M14 cbg_M14 cbd_M14 cbs_M14 cdg_M14 cdd_M14 cds_M14 csg_M14 csd_M14 css_M14 cgb_M14 cdb_M14 csb_M14 cbb_M14 capbd_M14 capbs_M14 gmbs_M15 gm_M15 gds_M15 vdsat_M15 vth_M15 id_M15 ibd_M15 ibs_M15 gbd_M15 gbs_M15 isub_M15 igidl_M15 igisl_M15 igs_M15 igd_M15 igb_M15 igcs_M15 vbs_M15 vgs_M15 vds_M15 cgg_M15 cgs_M15 cgd_M15 cbg_M15 cbd_M15 cbs_M15 cdg_M15 cdd_M15 cds_M15 csg_M15 csd_M15 css_M15 cgb_M15 cdb_M15 csb_M15 cbb_M15 capbd_M15 capbs_M15 gmbs_M16 gm_M16 gds_M16 vdsat_M16 vth_M16 id_M16 ibd_M16 ibs_M16 gbd_M16 gbs_M16 isub_M16 igidl_M16 igisl_M16 igs_M16 igd_M16 igb_M16 igcs_M16 vbs_M16 vgs_M16 vds_M16 cgg_M16 cgs_M16 cgd_M16 cbg_M16 cbd_M16 cbs_M16 cdg_M16 cdd_M16 cds_M16 csg_M16 csd_M16 css_M16 cgb_M16 cdb_M16 csb_M16 cbb_M16 capbd_M16 capbs_M16 gmbs_M17 gm_M17 gds_M17 vdsat_M17 vth_M17 id_M17 ibd_M17 ibs_M17 gbd_M17 gbs_M17 isub_M17 igidl_M17 igisl_M17 igs_M17 igd_M17 igb_M17 igcs_M17 vbs_M17 vgs_M17 vds_M17 cgg_M17 cgs_M17 cgd_M17 cbg_M17 cbd_M17 cbs_M17 cdg_M17 cdd_M17 cds_M17 csg_M17 csd_M17 css_M17 cgb_M17 cdb_M17 csb_M17 cbb_M17 capbd_M17 capbs_M17 gmbs_M18 gm_M18 gds_M18 vdsat_M18 vth_M18 id_M18 ibd_M18 ibs_M18 gbd_M18 gbs_M18 isub_M18 igidl_M18 igisl_M18 igs_M18 igd_M18 igb_M18 igcs_M18 vbs_M18 vgs_M18 vds_M18 cgg_M18 cgs_M18 cgd_M18 cbg_M18 cbd_M18 cbs_M18 cdg_M18 cdd_M18 cds_M18 csg_M18 csd_M18 css_M18 cgb_M18 cdb_M18 csb_M18 cbb_M18 capbd_M18 capbs_M18 gmbs_M19 gm_M19 gds_M19 vdsat_M19 vth_M19 id_M19 ibd_M19 ibs_M19 gbd_M19 gbs_M19 isub_M19 igidl_M19 igisl_M19 igs_M19 igd_M19 igb_M19 igcs_M19 vbs_M19 vgs_M19 vds_M19 cgg_M19 cgs_M19 cgd_M19 cbg_M19 cbd_M19 cbs_M19 cdg_M19 cdd_M19 cds_M19 csg_M19 csd_M19 css_M19 cgb_M19 cdb_M19 csb_M19 cbb_M19 capbd_M19 capbs_M19 gmbs_M20 gm_M20 gds_M20 vdsat_M20 vth_M20 id_M20 ibd_M20 ibs_M20 gbd_M20 gbs_M20 isub_M20 igidl_M20 igisl_M20 igs_M20 igd_M20 igb_M20 igcs_M20 vbs_M20 vgs_M20 vds_M20 cgg_M20 cgs_M20 cgd_M20 cbg_M20 cbd_M20 cbs_M20 cdg_M20 cdd_M20 cds_M20 csg_M20 csd_M20 css_M20 cgb_M20 cdb_M20 csb_M20 cbb_M20 capbd_M20 capbs_M20 gmbs_M21 gm_M21 gds_M21 vdsat_M21 vth_M21 id_M21 ibd_M21 ibs_M21 gbd_M21 gbs_M21 isub_M21 igidl_M21 igisl_M21 igs_M21 igd_M21 igb_M21 igcs_M21 vbs_M21 vgs_M21 vds_M21 cgg_M21 cgs_M21 cgd_M21 cbg_M21 cbd_M21 cbs_M21 cdg_M21 cdd_M21 cds_M21 csg_M21 csd_M21 css_M21 cgb_M21 cdb_M21 csb_M21 cbb_M21 capbd_M21 capbs_M21 gmbs_M22 gm_M22 gds_M22 vdsat_M22 vth_M22 id_M22 ibd_M22 ibs_M22 gbd_M22 gbs_M22 isub_M22 igidl_M22 igisl_M22 igs_M22 igd_M22 igb_M22 igcs_M22 vbs_M22 vgs_M22 vds_M22 cgg_M22 cgs_M22 cgd_M22 cbg_M22 cbd_M22 cbs_M22 cdg_M22 cdd_M22 cds_M22 csg_M22 csd_M22 css_M22 cgb_M22 cdb_M22 csb_M22 cbb_M22 capbd_M22 capbs_M22 gmbs_M23 gm_M23 gds_M23 vdsat_M23 vth_M23 id_M23 ibd_M23 ibs_M23 gbd_M23 gbs_M23 isub_M23 igidl_M23 igisl_M23 igs_M23 igd_M23 igb_M23 igcs_M23 vbs_M23 vgs_M23 vds_M23 cgg_M23 cgs_M23 cgd_M23 cbg_M23 cbd_M23 cbs_M23 cdg_M23 cdd_M23 cds_M23 csg_M23 csd_M23 css_M23 cgb_M23 cdb_M23 csb_M23 cbb_M23 capbd_M23 capbs_M23 dc_Ib acmag_Ib acphase_Ib acreal_Ib acimag_Ib v_Ib p_Ib current_Ib capacitance_C0 cap_C0 c_C0 ic_C0 temp_C0 dtemp_C0 w_C0 l_C0 m_C0 scale_C0 i_C0 p_C0 sens_dc_C0 sens_real_C0 sens_imag_C0 sens_mag_C0 sens_ph_C0 sens_cplx_C0 capacitance_C1 cap_C1 c_C1 ic_C1 temp_C1 dtemp_C1 w_C1 l_C1 m_C1 scale_C1 i_C1 p_C1 sens_dc_C1 sens_real_C1 sens_imag_C1 sens_mag_C1 sens_ph_C1 sens_cplx_C1 

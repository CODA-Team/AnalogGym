.param MOSFET_0_8_W_BIASCM_PMOS=8.401687951475711 MOSFET_0_8_L_BIASCM_PMOS=1.8753550832847838 MOSFET_0_8_M_BIASCM_PMOS=19
.param MOSFET_8_2_W_gm1_PMOS=1.3222527842051277 MOSFET_8_2_L_gm1_PMOS=2.6270257845071705 MOSFET_8_2_M_gm1_PMOS=37
.param MOSFET_10_1_W_gm2_PMOS=1.710426467813417 MOSFET_10_1_L_gm2_PMOS=1.8154329552478603 MOSFET_10_1_M_gm2_PMOS=4
.param MOSFET_11_1_W_gmf2_PMOS=3.578620867067523 MOSFET_11_1_L_gmf2_PMOS=3.581661795317242 MOSFET_11_1_M_gmf2_PMOS=347
.param MOSFET_17_7_W_BIASCM_NMOS=1.4611546975877676 MOSFET_17_7_L_BIASCM_NMOS=0.9503514834662219 MOSFET_17_7_M_BIASCM_NMOS=4
.param MOSFET_21_2_W_LOAD2_NMOS=5.923108683557338 MOSFET_21_2_L_LOAD2_NMOS=1.3873797864025055 MOSFET_21_2_M_LOAD2_NMOS=42
.param MOSFET_23_1_W_gm3_NMOS=1.2341762562343073 MOSFET_23_1_L_gm3_NMOS=2.38420311655875 MOSFET_23_1_M_gm3_NMOS=9
.param CURRENT_0_BIAS=5.245106465782526e-06
.param M_C0=21
.param M_C1=8

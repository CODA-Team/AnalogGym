Test LDO ACDC

*.OPTIONS RELTOL=.0001
***************************************
* Step 1: Replace circuit netlist here.
*************************************** 
.include ../spice_netlist/LDO_netlist.txt

.param mc_mm_switch=0
.param mc_pr_switch=0

.include ../mosfet_model/sky130_pdk/libs.tech/ngspice/corners/tt.spice
.include ../mosfet_model/sky130_pdk/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ../mosfet_model/sky130_pdk/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ../mosfet_model/sky130_pdk/libs.tech/ngspice/corners/tt/specialized_cells.spice

***************************************
* Step 2: Replace circuit param.  here.
***************************************
.include ../design_variables/LDO_variables.txt
.PARAM supply_voltage = 1.8
.PARAM Vref = 0.4
.PARAM PARAM_ILOAD =55m 

V1 vdd 0 'supply_voltage'
V2 vss 0 0 

Vindc vref_in 0 'Vref'
Vin signal_in 0 dc 'Vref' ac 1 sin('Vref' 100m 500)

* Circuit List:
* Basic_LDO

* XLDO gnda vdda vinn vout vfb vinp Ib
*        |  |     |     |   |    |   |
*        |  |     |     |   |    |   bias current
*        |  |     |     |   |    Non-inverting input 
*        |  |     |     |   Feedback voltage 
*        |  |     |     |   
*        |  |     |     Output
*        |  |     Inverting Input
*        |  Positive Supply
*         Negative Supply 

***************************************
* Step 3: Replace circuit name below.
* e.g. Basic_LDO -> DFCFC_LDO
*************************************** 
*    ADM TB   
x1 vss vdd vref_in vout1 vfb1 vinp1 Ib Basic_LDO
Ib Ib 0 DC='current_0_bias'
Lfb vinp1 vfb1 1T
Cfb vinp1 signal_in 1T
XCL vout1 0 sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=M_CL m=M_CL
Iload1 vout1 0 'PARAM_ILOAD'

* PSRR   TB   
VVDDApsrr vddpsrr 0 'supply_voltage'  AC=1
Ib2 Ib2 0 DC='current_0_bias'
XCL2 ppsr1 0 sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=M_CL m=M_CL
x2 vss vddpsrr vref_in ppsr1 vfb2 vfb2 Ib2 Basic_LDO
Iload2 ppsr1 0 'PARAM_ILOAD'

* DC ALL  TB  
VVDDdc VDDdc 0 'supply_voltage' 
Ib3 Ib3 0 DC='current_0_bias'
XCL3 vout6 0 sky130_fd_pr__cap_mim_m3_1 W=30 L=30 MF=M_CL m=M_CL
x3 vss vdddc vref_in vout6 vfb3 vfb3 Ib3 Basic_LDO
Iload3 vout6 0 'PARAM_ILOAD'

.control
* save all voltage and current
save all
.options savecurrents 
set filetype=ascii
set units=degrees

* LNR at maxload
alter Iload3 dc=55m
dc VVDDdc 1.62 1.98 0.01
meas dc maxval1 MAX V(vout6) from=1.62 to=1.98
meas dc minval1 MIN V(vout6) from=1.62 to=1.98
meas dc avgval1 AVG V(vout6) from=1.62 to=1.98
meas dc ppavl1  PP V(vout6) from=1.62 to=1.98
let LNR1 = ppavl1/avgval1/0.36
print LNR1
plot v(vout6)
wrdata LDO_TB_ACDC_LNR_maxload LNR1

* LNR at minload
alter Iload3 dc=5m
dc VVDDdc 1.62 1.98 0.01
meas dc maxval2 MAX V(vout6) from=1.62 to=1.98
meas dc minval2 MIN V(vout6) from=1.62 to=1.98
meas dc avgval2 AVG V(vout6) from=1.62 to=1.98
meas dc ppavl2  PP V(vout6) from=1.62 to=1.98
let LNR2 = ppavl2/avgval2/0.36
print LNR2
plot v(vout6)
wrdata LDO_TB_ACDC_LNR_minload LNR2

dc Iload3 5m 55m 0.1m
* LR meas   
meas dc maxval MAX V(vout6) from=5m to=55m
meas dc minval MIN V(vout6) from=5m to=55m
meas dc avgval AVG V(vout6) from=5m to=55m
meas dc ppavl  PP V(vout6) from=5m to=55m
let LR = ppavl/avgval/50m
print LR
* Power meas at maxload
meas dc Ivdd1 FIND I(VVDDDC) AT=55m
let Power1 = -1*Ivdd1*1.8
print Power1
* Power meas at minload
meas dc Ivdd2 FIND I(VVDDDC) AT=5m
let Power2 = -1*Ivdd2*1.8
print Power2
*   Vos.meas at maxload
meas dc vout_x FIND V(vout6) AT=55m
let vos1 = vout_x-4*0.4
print vos1
*   Vos.meas at minload
meas dc vout_y FIND V(vout6) AT=5m
let vos2 = vout_y-4*0.4
print vos2
plot v(vout6)
wrdata LDO_TB_ACDC_LR_Power_vos LR Power1 Power2 vos1 vos2 

* Loop test at maxload
alter Iload1 dc=55m
ac dec 10 0.1 1G
meas ac DCPSRp1 find vdb(ppsr1) at = 0.1
meas ac dcgain1 find vdb(vout1) at = 0.1
meas ac gain_bandwidth_product1 when vdb(vout1)=0
meas ac phase_margin1 find vp(vout1) when vdb(vout1)=0
plot vdb(vout1) vdb(ppsr1) vp(vout1)
wrdata LDO_TB_ACDC_PSRR_dcgain_maxload DCPSRp1 dcgain1
wrdata LDO_TB_ACDC_GBW_PM_maxload gain_bandwidth_product1 phase_margin1

* Loop test at minload
alter Iload1 dc=5m
ac dec 10 0.1 1G
meas ac DCPSRp2 find vdb(ppsr1) at = 0.1
meas ac dcgain2 find vdb(vout1) at = 0.1
meas ac gain_bandwidth_product2 when vdb(vout1)=0
meas ac phase_margin2 find vp(vout1) when vdb(vout1)=0
plot vdb(vout1) vdb(ppsr1) vp(vout1)
wrdata LDO_TB_ACDC_PSRR_dcgain_minload DCPSRp2 dcgain2
wrdata LDO_TB_ACDC_GBW_PM_minload gain_bandwidth_product2 phase_margin2

.endc

.end

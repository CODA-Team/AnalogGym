Test OpAmp Tran

*.OPTIONS RELTOL=.0001
***************************************
* Step 1: Replace circuit netlist here.
*************************************** 
*.include ./netlist/NMCNR_Pin_3_HSPICE.txt
.include ./netlist/NMCNR_Pin_3_HSPICE_130.txt
*.include ./netlist/NMCF_Pin_3_HSPICE.txt
*.include ./netlist/DFCFC1_Pin_3_HSPICE.txt
*.include ./netlist/DFCFC2_Pin_3_HSPICE.txt


*.include ./mosfet_model/modelcard.nmos
*.include ./mosfet_model/modelcard.pmos

.param mc_mm_switch=0
.param mc_pr_switch=0

.include ./mosfet_model/sky130_pdk/libs.tech/ngspice/corners/tt.spice
*.include.\mosfet_model\sky130_pdk\libs.tech\ngspice\r+c\res_typical__cap_typical.spice
*.include.\mosfet_model\sky130_pdk\libs.tech\ngspice\r+c\res_typical__cap_typical__lin.spice
*.include.\mosfet_model\sky130_pdk\libs.tech\ngspice\corners\tt\specialized_cells.spice


.PARAM supply_voltage = 1.8
.PARAM VCM_ratio = 0.4
.PARAM PARAM_CLOAD =100.00p 
.PARAM val0 = 3.000000e-01
.PARAM val1 = 5.000000e-01
.PARAM GBW_ideal = 5e4
.PARAM STEP_TIME = '10/GBW_ideal'
.PARAM TRAN_SIM_TIME = '20/GBW_ideal + 1e-6'


***************************************
* Step 2: Replace circuit param.  here.
*************************************** 
*NMCNR 
*.PARAM RESISTOR_0=0.5k MOSFET_10_1_L_gm2_PMOS=1u MOSFET_10_1_M_gm2_PMOS=38  
*+ MOSFET_10_1_W_gm2_PMOS=0.5u MOSFET_23_1_L_gm3_NMOS=1u MOSFET_23_1_M_gm3_NMOS=40  
*+ MOSFET_23_1_W_gm3_NMOS=0.5u MOSFET_8_2_L_gm1_PMOS=1u MOSFET_8_2_M_gm1_PMOS=37  
*+ MOSFET_8_2_W_gm1_PMOS=0.5u MOSFET_0_8_L_BIASCM_PMOS=1u MOSFET_0_8_M_BIASCM_PMOS=40  
*+ MOSFET_0_8_W_BIASCM_PMOS=0.5u MOSFET_17_7_L_BIASCM_NMOS=1u MOSFET_17_7_M_BIASCM_NMOS=10  
*+ MOSFET_17_7_W_BIASCM_NMOS=0.5u MOSFET_21_2_L_LOAD2_NMOS=1u MOSFET_21_2_M_LOAD2_NMOS=25  
*+ MOSFET_21_2_W_LOAD2_NMOS=0.411u CAPACITOR_0=63p CAPACITOR_1=25p  
*+ CURRENT_0_BIAS=5u

.PARAM RESISTOR_0=0.5k MOSFET_10_1_L_gm2_PMOS=0.5 
 +MOSFET_10_1_M_gm2_PMOS=193.0 MOSFET_10_1_W_gm2_PMOS=1.01 
 +MOSFET_23_1_L_gm3_NMOS=0.5 MOSFET_23_1_M_gm3_NMOS=200.0 
 +MOSFET_23_1_W_gm3_NMOS=1.0 MOSFET_8_2_L_gm1_PMOS=0.5
 +MOSFET_8_2_M_gm1_PMOS=183.0 MOSFET_8_2_W_gm1_PMOS=1.0
 +MOSFET_0_8_L_BIASCM_PMOS=0.5 MOSFET_0_8_M_BIASCM_PMOS=200.0 
 +MOSFET_0_8_W_BIASCM_PMOS=1.0 MOSFET_17_7_L_BIASCM_NMOS=0.5 
 +MOSFET_17_7_M_BIASCM_NMOS=1.0 MOSFET_17_7_W_BIASCM_NMOS=1.01 
 +MOSFET_21_2_L_LOAD2_NMOS=1.0 MOSFET_21_2_M_LOAD2_NMOS=125.0 
 +MOSFET_21_2_W_LOAD2_NMOS=0.645 CAPACITOR_0=63.0p CAPACITOR_1=25.0p 
 +CURRENT_0_BIAS=5.0u


*NMCF
*.PARAM MOSFET_10_1_L_gm2_PMOS=1u MOSFET_10_1_M_gm2_PMOS=13 MOSFET_10_1_W_gm2_PMOS=0.99u  
*+ MOSFET_11_1_L_gmf2_PMOS=1u MOSFET_11_1_M_gmf2_PMOS=333 MOSFET_11_1_W_gmf2_PMOS=1u  
*+ MOSFET_23_1_L_gm3_NMOS=1u MOSFET_23_1_M_gm3_NMOS=47 MOSFET_23_1_W_gm3_NMOS=1u  
*+ MOSFET_8_2_L_gm1_PMOS=1u MOSFET_8_2_M_gm1_PMOS=13 MOSFET_8_2_W_gm1_PMOS=0.99u  
*+ MOSFET_0_8_L_BIASCM_PMOS=1u MOSFET_0_8_M_BIASCM_PMOS=24 MOSFET_0_8_W_BIASCM_PMOS=1u  
*+ MOSFET_17_7_L_BIASCM_NMOS=1u MOSFET_17_7_M_BIASCM_NMOS=11 MOSFET_17_7_W_BIASCM_NMOS=0.97u  
*+ MOSFET_21_2_L_LOAD2_NMOS=1u MOSFET_21_2_M_LOAD2_NMOS=1 MOSFET_21_2_W_LOAD2_NMOS=2.14667u  
*+ CAPACITOR_0=7.14p CAPACITOR_1=11.3p CURRENT_0_BIAS=1u  

*DFCFC1 
*.PARAM MOSFET_0_8_L_BIASCM_PMOS=1u MOSFET_0_8_M_BIASCM_PMOS=45 MOSFET_0_8_W_BIASCM_PMOS=1u  
*+ MOSFET_11_1_L_gm2_PMOS=1u MOSFET_11_1_M_gm2_PMOS=14 MOSFET_11_1_W_gm2_PMOS=0.99u  
*+ MOSFET_12_1_L_gmf2_PMOS=1u MOSFET_12_1_M_gmf2_PMOS=240 MOSFET_12_1_W_gmf2_PMOS=1u  
*+ MOSFET_17_7_L_BIASCM_NMOS=1u MOSFET_17_7_M_BIASCM_NMOS=40 MOSFET_17_7_W_BIASCM_NMOS=0.98u  
*+ MOSFET_18_7_L_BIASCM_NMOS=1u MOSFET_18_7_M_BIASCM_NMOS=8 MOSFET_18_7_W_BIASCM_NMOS=0.99u  
*+ MOSFET_22_2_L_LOAD2_NMOS=1u MOSFET_22_2_M_LOAD2_NMOS=5 MOSFET_22_2_W_LOAD2_NMOS=0.88u  
*+ MOSFET_24_1_L_gm4_NMOS=1u MOSFET_24_1_M_gm4_NMOS=1 MOSFET_24_1_W_gm4_NMOS=0.942u  
*+ MOSFET_25_1_L_gm3_NMOS=1u MOSFET_25_1_M_gm3_NMOS=16 MOSFET_25_1_W_gm3_NMOS=1u  
*+ MOSFET_9_2_L_gm1_PMOS=1u MOSFET_9_2_M_gm1_PMOS=17 MOSFET_9_2_W_gm1_PMOS=0.99u  
*+ CAPACITOR_0=3.85p CAPACITOR_1=0.5p CURRENT_0_BIAS=5u  

*DFCFC2
*.PARAM MOSFET_0_8_L_BIASCM_PMOS=1u MOSFET_0_8_M_BIASCM_PMOS=10 MOSFET_0_8_W_BIASCM_PMOS=0.98u  
*+ MOSFET_10_1_L_gm4_PMOS=1u MOSFET_10_1_M_gm4_PMOS=1 MOSFET_10_1_W_gm4_PMOS=2.352u  
*+ MOSFET_11_1_L_gm2_PMOS=1u MOSFET_11_1_M_gm2_PMOS=1 MOSFET_11_1_W_gm2_PMOS=0.792u  
*+ MOSFET_12_1_L_gmf2_PMOS=1u MOSFET_12_1_M_gmf2_PMOS=17 MOSFET_12_1_W_gmf2_PMOS=1u  
*+ MOSFET_18_7_L_BIASCM_NMOS=1u MOSFET_18_7_M_BIASCM_NMOS=6 MOSFET_18_7_W_BIASCM_NMOS=0.99u  
*+ MOSFET_23_2_L_LOAD2_NMOS=1u MOSFET_23_2_M_LOAD2_NMOS=1 MOSFET_23_2_W_LOAD2_NMOS=4.158u  
*+ MOSFET_25_1_L_gm3_NMOS=1u MOSFET_25_1_M_gm3_NMOS=6 MOSFET_25_1_W_gm3_NMOS=0.98u  
*+ MOSFET_8_2_L_gm1_PMOS=1u MOSFET_8_2_M_gm1_PMOS=7 MOSFET_8_2_W_gm1_PMOS=0.98u  
*+ CAPACITOR_0=3.85p CAPACITOR_1=0.5p CURRENT_0_BIAS=2.3u  


V1 vdd 0 'supply_voltage'
V2 vss 0 0 

* Circuit List:
* Leung_NMCNR_Pin_3
* Leung_NMCF_Pin_3
* Leung_DFCFC1_Pin_3
* Leung_DFCFC2_Pin_3

* XOP gnda vdda vinn vinp vout
*        |  |     |     |   |
*        |  |     |     |   Output
*        |  |     |     Non-inverting Input
*        |  |      Inverting Input
*        |  Positive Supply
*        Negative Supply 

***************************************
* Step 3: Replace circuit name below.
* e.g. Leung_NMCNR_Pin_3 -> Leung_NMCF_Pin_3
*************************************** 
*Transient  TB  
VVISR visr 0 pulse('val0' 'val1' 1u 1p 1p '1*STEP_TIME' 1)
xop6 vss vdd vout3 visr vout3 Leung_NMCNR_Pin_3
CLoad6 vout3 0 'PARAM_CLOAD'

.meas tran t_rise_edge when v(vout3)=0.4 rise=1
.meas tran t_rise param='t_rise_edge-1u'
.meas tran sr_rise param='0.1/t_rise'

.meas tran t_fall_edge when v(vout3)=0.4 fall=1
.meas tran t_fall param='t_fall_edge-1u-STEP_TIME'
.meas tran sr_fall param='0.1/t_fall'

.control

tran 1u 4.01e-4
plot v(visr) v(vout3)
write tran.dat v(vout3)
.endc

.end

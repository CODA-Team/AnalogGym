Test LDO Tran

*.OPTIONS RELTOL=.0001
***************************************
* Step 1: Replace circuit netlist here.
*************************************** 
.include ./ldo_spice_netlist/LDO_1.txt
.include ./ldo_spice_parameter/LDO_1.txt

.param mc_mm_switch=0
.param mc_pr_switch=0

.include ./mosfet_model/sky130_pdk/libs.tech/ngspice/corners/tt.spice
*.include.\mosfet_model\sky130_pdk\libs.tech\ngspice\r+c\res_typical__cap_typical.spice
*.include.\mosfet_model\sky130_pdk\libs.tech\ngspice\r+c\res_typical__cap_typical__lin.spice
*.include.\mosfet_model\sky130_pdk\libs.tech\ngspice\corners\tt\specialized_cells.spice

.PARAM supply_voltage = 1.8
.PARAM Vref = 0.4
.PARAM PARAM_CLOAD =100.00p 
.PARAM PARAM_ILOAD =10n 
.PARAM val0 = 1n
.PARAM val1 = 5m
.PARAM GBW_ideal = 5e4
.PARAM STEP_TIME = '10/GBW_ideal'


V1 vdd 0 'supply_voltage'
V2 vss 0 0 

Vindc vref_in 0 'Vref'

* Circuit List:
* Basic_LDO


* XLDO gnda vdda vinn vout vddp vfb vinp
*        |  |     |     |   |    |   |
*        |  |     |     |   |    |   Non-inverting input
*        |  |     |     |   |    Feedback voltage 
*        |  |     |     |   Supply of the Power transistor
*        |  |     |     Output
*        |  |      Inverting Input
*        |  Positive Supply
*        Negative Supply 

***************************************
* Step 3: Replace circuit name below.
* e.g. Basic_LDO -> DFCFC_LDO
*************************************** 
*   Tran TB   
Xldo1 vss vdd vref_in vout1 vdd vfb1 vfb1 Basic_LDO
Cload1 vout1 0 'PARAM_CLOAD'
Iload1 vout1 0 pulse('val0' 'val1' 1u 1p 1p '1*STEP_TIME' 1)

.meas tran v_min MIN v(vout1) from=900n to='900n+STEP_TIME'
.meas tran v_max MAX v(vout1) from='900n+STEP_TIME' to=1m
.meas tran v_undershoot param='4*vref - v_min'
.meas tran v_overshoot param='v_max - 4*vref'

*   Voltage Regulation meas 
.measure dc maxval MAX V(vout1) from='0.9*Vref*4' to='1.1*Vref*4'
.measure dc minval MIN V(vout1) from='0.9*Vref*4' to='1.1*Vref*4'
.measure dc avgval AVG V(vout1) from='0.9*Vref*4' to='1.1*Vref*4'
.measure dc ppavl  PP V(vout1) from='0.9*Vref*4' to='1.1*Vref*4'
.measure dc VR param='ppavl/avgval/0.8/Vref'

.control

tran 1u 1m
dc v1 0 2 0.1
plot v(vout1)
write tran.dat v(vout1)

.endc

.end
